----------------------------------------------------------------------------
--
--  Copyright (c) 2013, Tom Hunter
--
--  Project     : CDC 6612 display controller
--  File        : char_rom.vhd
--  Description : Character ROM for DD60 console glyphs.
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License version 3 as
--  published by the Free Software Foundation.
--  
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License version 3 for more details.
--  
--  You should have received a copy of the GNU General Public License
--  version 3 along with this program in file "license-gpl-3.0.txt".
--  If not, see <http://www.gnu.org/licenses/gpl-3.0.txt>.
--
----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use work.controller.all;

entity char_rom is 
port
(
  clk_10mhz     : in std_logic;
  char          : in integer range 0 to (char_rom_chars - 1);
  row           : in integer range 0 to (char_rom_rows - 1);
  data          : out std_logic_vector((char_rom_bits - 1) downto 0)
);

end;

architecture behavior of char_rom is
type rom_type is array (0 to (char_rom_words - 1)) of std_logic_vector ((char_rom_bits - 1) downto 0);
signal read_data : std_logic_vector ((char_rom_bits - 1) downto 0);
signal rom : rom_type:=
(
  -- ' ' (00)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'A' (01)
  "00000", -- 76 
  "00001", -- 00 
  "01100", -- 01 
  "01100", -- 02 
  "01100", -- 03 
  "11000", -- 04 
  "01100", -- 05 
  "01100", -- 06 
  "01100", -- 07 
  "11110", -- 10 
  "01101", -- 11 
  "00001", -- 12 
  "00010", -- 13 
  "00010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'B' (02)
  "00001", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11000", -- 03 
  "00010", -- 04 
  "00010", -- 05 
  "10010", -- 06 
  "10110", -- 07 
  "10010", -- 10 
  "00010", -- 11 
  "00010", -- 12 
  "00110", -- 13 
  "00011", -- 14 
  "00011", -- 15 
  "10010", -- 16 
  "10110", -- 17 
  "10010", -- 20 
  "00010", -- 21 
  "00010", -- 22 
  "00000", -- 23 
  "00001", -- 24 
  "00000", -- 25 

  -- 'C' (03)
  "01010", -- 76 
  "01010", -- 00 
  "10010", -- 01 
  "00000", -- 02 
  "00111", -- 03 
  "10010", -- 04 
  "11010", -- 05 
  "10010", -- 06 
  "01110", -- 07 
  "01000", -- 10 
  "10010", -- 11 
  "11010", -- 12 
  "10010", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'D' (04)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11000", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "10010", -- 07 
  "01110", -- 10 
  "01000", -- 11 
  "10010", -- 12 
  "00010", -- 13 
  "00010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'E' (05)
  "00001", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11000", -- 03 
  "00010", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "00111", -- 07 
  "01010", -- 10 
  "00000", -- 11 
  "00011", -- 12 
  "00010", -- 13 
  "00110", -- 14 
  "01001", -- 15 
  "01000", -- 16 
  "00001", -- 17 
  "00010", -- 20 
  "00010", -- 21 
  "00010", -- 22 
  "00000", -- 23 
  "00001", -- 24 
  "00000", -- 25 

  -- 'F' (06)
  "00001", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11000", -- 03 
  "00010", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "00111", -- 07 
  "01010", -- 10 
  "10000", -- 11 
  "00000", -- 12 
  "00011", -- 13 
  "00010", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'G' (07)
  "10010", -- 76 
  "01010", -- 00 
  "00000", -- 01 
  "00001", -- 02 
  "00010", -- 03 
  "11110", -- 04 
  "01000", -- 05 
  "10010", -- 06 
  "11010", -- 07 
  "10010", -- 10 
  "01110", -- 11 
  "01000", -- 12 
  "10010", -- 13 
  "11010", -- 14 
  "10010", -- 15 
  "00000", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'H' (10)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11001", -- 04 
  "01000", -- 05 
  "10001", -- 06 
  "00000", -- 07 
  "00010", -- 10 
  "00010", -- 11 
  "00010", -- 12 
  "00000", -- 13 
  "01001", -- 14 
  "10000", -- 15 
  "11001", -- 16 
  "01000", -- 17 
  "01000", -- 20 
  "01000", -- 21 
  "00000", -- 22 
  "00001", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'I' (11)
  "00010", -- 76 
  "00100", -- 00 
  "00001", -- 01 
  "00000", -- 02 
  "01000", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "00001", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'J' (12)
  "01000", -- 76 
  "11001", -- 00 
  "01010", -- 01 
  "11010", -- 02 
  "01010", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "00001", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'K' (13)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11001", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "00011", -- 07 
  "00110", -- 10 
  "10010", -- 11 
  "10010", -- 12 
  "10010", -- 13 
  "00110", -- 14 
  "10010", -- 15 
  "10010", -- 16 
  "10010", -- 17 
  "00000", -- 20 
  "00001", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'L' (14)
  "00000", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11001", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "01000", -- 06 
  "00000", -- 07 
  "00010", -- 10 
  "00010", -- 11 
  "00010", -- 12 
  "00000", -- 13 
  "00001", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'M' (15)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11000", -- 04 
  "01010", -- 05 
  "10100", -- 06 
  "11000", -- 07 
  "01010", -- 10 
  "10100", -- 11 
  "11000", -- 12 
  "01000", -- 13 
  "01000", -- 14 
  "01000", -- 15 
  "00000", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'N' (16)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11000", -- 04 
  "01010", -- 05 
  "01010", -- 06 
  "01010", -- 07 
  "11000", -- 10 
  "01000", -- 11 
  "01000", -- 12 
  "01000", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'O' (17)
  "01000", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "01000", -- 02 
  "01010", -- 03 
  "11010", -- 04 
  "01010", -- 05 
  "01110", -- 06 
  "01010", -- 07 
  "11010", -- 10 
  "01010", -- 11 
  "00001", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'P' (20)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11000", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "10010", -- 07 
  "10110", -- 10 
  "10010", -- 11 
  "00010", -- 12 
  "00010", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'Q' (21)
  "00010", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "00010", -- 02 
  "01010", -- 03 
  "01110", -- 04 
  "01010", -- 05 
  "11010", -- 06 
  "01010", -- 07 
  "01110", -- 10 
  "01010", -- 11 
  "11001", -- 12 
  "01010", -- 13 
  "11000", -- 14 
  "00001", -- 15 
  "01010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'R' (22)
  "00000", -- 76 
  "00001", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "11000", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "10010", -- 07 
  "10110", -- 10 
  "10010", -- 11 
  "00010", -- 12 
  "00010", -- 13 
  "00110", -- 14 
  "10010", -- 15 
  "10010", -- 16 
  "10010", -- 17 
  "00000", -- 20 
  "00001", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'S' (23)
  "10000", -- 76 
  "00000", -- 00 
  "11001", -- 01 
  "10010", -- 02 
  "11010", -- 03 
  "10010", -- 04 
  "10110", -- 05 
  "10010", -- 06 
  "00010", -- 07 
  "10010", -- 10 
  "10110", -- 11 
  "10010", -- 12 
  "11010", -- 13 
  "10010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'T' (24)
  "00010", -- 76 
  "00100", -- 00 
  "00000", -- 01 
  "00001", -- 02 
  "01000", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "00001", -- 06 
  "00010", -- 07 
  "00100", -- 10 
  "00111", -- 11 
  "00010", -- 12 
  "00010", -- 13 
  "00010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'U' (25)
  "00000", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11001", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "01100", -- 06 
  "11010", -- 07 
  "00010", -- 10 
  "01100", -- 11 
  "01000", -- 12 
  "01000", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'V' (26)
  "00000", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11001", -- 03 
  "01100", -- 04 
  "01100", -- 05 
  "01100", -- 06 
  "11000", -- 07 
  "01100", -- 10 
  "01100", -- 11 
  "01100", -- 12 
  "00000", -- 13 
  "00001", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'W' (27)
  "00000", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "01000", -- 02 
  "11001", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "01000", -- 06 
  "11000", -- 07 
  "01010", -- 10 
  "10100", -- 11 
  "11000", -- 12 
  "01010", -- 13 
  "10100", -- 14 
  "11000", -- 15 
  "01000", -- 16 
  "01000", -- 17 
  "01000", -- 20 
  "00000", -- 21 
  "00001", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'X' (30)
  "00000", -- 76 
  "00001", -- 00 
  "01010", -- 01 
  "01010", -- 02 
  "01010", -- 03 
  "11111", -- 04 
  "01000", -- 05 
  "01000", -- 06 
  "01000", -- 07 
  "11001", -- 10 
  "01010", -- 11 
  "01010", -- 12 
  "01010", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'Y' (31)
  "00010", -- 76 
  "00100", -- 00 
  "00000", -- 01 
  "00001", -- 02 
  "01000", -- 03 
  "10000", -- 04 
  "00001", -- 05 
  "01010", -- 06 
  "10100", -- 07 
  "11111", -- 10 
  "01010", -- 11 
  "10100", -- 12 
  "11000", -- 13 
  "01010", -- 14 
  "10100", -- 15 
  "00000", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- 'Z' (32)
  "01000", -- 76 
  "01000", -- 00 
  "01000", -- 01 
  "00000", -- 02 
  "11001", -- 03 
  "00010", -- 04 
  "00010", -- 05 
  "00010", -- 06 
  "00110", -- 07 
  "01010", -- 10 
  "01010", -- 11 
  "01010", -- 12 
  "00110", -- 13 
  "00010", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '0' (33)
  "10000", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "01000", -- 02 
  "01000", -- 03 
  "10100", -- 04 
  "11010", -- 05 
  "00010", -- 06 
  "10100", -- 07 
  "01110", -- 10 
  "01000", -- 11 
  "10100", -- 12 
  "11010", -- 13 
  "00010", -- 14 
  "10100", -- 15 
  "00000", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '1' (34)
  "00010", -- 76 
  "00100", -- 00 
  "00000", -- 01 
  "00111", -- 02 
  "01000", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "11000", -- 06 
  "10010", -- 07 
  "00000", -- 10 
  "00001", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '2' (35)
  "01000", -- 76 
  "01000", -- 00 
  "10000", -- 01 
  "00000", -- 02 
  "00001", -- 03 
  "10010", -- 04 
  "11010", -- 05 
  "10010", -- 06 
  "10110", -- 07 
  "10010", -- 10 
  "10010", -- 11 
  "01010", -- 12 
  "00110", -- 13 
  "00010", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '3' (36)
  "10000", -- 76 
  "00000", -- 00 
  "11001", -- 01 
  "10010", -- 02 
  "11010", -- 03 
  "10010", -- 04 
  "01110", -- 05 
  "10010", -- 06 
  "00010", -- 07 
  "00110", -- 10 
  "10010", -- 11 
  "10010", -- 12 
  "00110", -- 13 
  "00010", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '4' (37)
  "00010", -- 76 
  "00010", -- 00 
  "00000", -- 01 
  "00111", -- 02 
  "01000", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "11000", -- 06 
  "01010", -- 07 
  "01010", -- 10 
  "00110", -- 11 
  "00010", -- 12 
  "00010", -- 13 
  "00010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '5' (40)
  "10000", -- 76 
  "00000", -- 00 
  "11001", -- 01 
  "10010", -- 02 
  "11010", -- 03 
  "10010", -- 04 
  "01110", -- 05 
  "10010", -- 06 
  "00010", -- 07 
  "00010", -- 10 
  "00000", -- 11 
  "01110", -- 12 
  "00000", -- 13 
  "00010", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '6' (41)
  "00000", -- 76 
  "01000", -- 00 
  "10000", -- 01 
  "00001", -- 02 
  "10010", -- 03 
  "11010", -- 04 
  "10010", -- 05 
  "01110", -- 06 
  "10010", -- 07 
  "11010", -- 10 
  "10010", -- 11 
  "01110", -- 12 
  "01000", -- 13 
  "10010", -- 14 
  "11010", -- 15 
  "10010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '7' (42)
  "00010", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "10000", -- 02 
  "01100", -- 03 
  "01010", -- 04 
  "10100", -- 05 
  "00110", -- 06 
  "00010", -- 07 
  "00010", -- 10 
  "00010", -- 11 
  "00001", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '8' (43)
  "10000", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "10000", -- 02 
  "10010", -- 03 
  "00010", -- 04 
  "10010", -- 05 
  "10110", -- 06 
  "10010", -- 07 
  "11010", -- 10 
  "10010", -- 11 
  "10110", -- 12 
  "10010", -- 13 
  "00010", -- 14 
  "10010", -- 15 
  "10110", -- 16 
  "10010", -- 17 
  "11010", -- 20 
  "10010", -- 21 
  "00000", -- 22 
  "00001", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '9' (44)
  "10000", -- 76 
  "00000", -- 00 
  "11001", -- 01 
  "10010", -- 02 
  "11010", -- 03 
  "10010", -- 04 
  "01110", -- 05 
  "01000", -- 06 
  "10010", -- 07 
  "11010", -- 10 
  "10010", -- 11 
  "01110", -- 12 
  "10010", -- 13 
  "11010", -- 14 
  "10010", -- 15 
  "00000", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '+' (45)
  "00010", -- 76 
  "00100", -- 00 
  "00000", -- 01 
  "00001", -- 02 
  "01000", -- 03 
  "01000", -- 04 
  "01000", -- 05 
  "11001", -- 06 
  "01010", -- 07 
  "10100", -- 10 
  "00111", -- 11 
  "00010", -- 12 
  "00010", -- 13 
  "00010", -- 14 
  "00000", -- 15 
  "00001", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '-' (46)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "01000", -- 07 
  "10000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00001", -- 13 
  "00010", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '*' (47)
  "10000", -- 76 
  "00100", -- 00 
  "00001", -- 01 
  "01010", -- 02 
  "01010", -- 03 
  "11111", -- 04 
  "01000", -- 05 
  "00001", -- 06 
  "00010", -- 07 
  "00010", -- 10 
  "11110", -- 11 
  "01001", -- 12 
  "11000", -- 13 
  "00001", -- 14 
  "01010", -- 15 
  "01010", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '/' (50)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00001", -- 14 
  "01010", -- 15 
  "01010", -- 16 
  "01010", -- 17 
  "00000", -- 20 
  "00001", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '(' (51)
  "00010", -- 76 
  "00010", -- 00 
  "00000", -- 01 
  "00111", -- 02 
  "10100", -- 03 
  "01110", -- 04 
  "01000", -- 05 
  "10100", -- 06 
  "00000", -- 07 
  "00001", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- ')' (52)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00010", -- 10 
  "00000", -- 11 
  "00001", -- 12 
  "10100", -- 13 
  "01110", -- 14 
  "01000", -- 15 
  "10100", -- 16 
  "00001", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- ' ' (53)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '=' (54)
  "01000", -- 76 
  "00000", -- 00 
  "00001", -- 01 
  "00010", -- 02 
  "00010", -- 03 
  "00010", -- 04 
  "00111", -- 05 
  "01000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00001", -- 14 
  "00010", -- 15 
  "00010", -- 16 
  "00010", -- 17 
  "00000", -- 20 
  "00001", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- ' ' (55)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00000", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00000", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- ',' (56)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00001", -- 14 
  "10100", -- 15 
  "11000", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000", -- 25 

  -- '.' (57)
  "00000", -- 76 
  "00000", -- 00 
  "00000", -- 01 
  "00000", -- 02 
  "00000", -- 03 
  "00000", -- 04 
  "00000", -- 05 
  "00000", -- 06 
  "00000", -- 07 
  "00000", -- 10 
  "00000", -- 11 
  "00000", -- 12 
  "00000", -- 13 
  "00000", -- 14 
  "00001", -- 15 
  "00000", -- 16 
  "00000", -- 17 
  "00001", -- 20 
  "00000", -- 21 
  "00000", -- 22 
  "00000", -- 23 
  "00000", -- 24 
  "00000"  -- 25 
);

begin

  read_data <= rom((char * char_rom_rows) + row) when char < char_rom_chars else "00000";

  read_row: process (clk_10mhz, char, row)
  begin
    if (rising_edge(clk_10mhz)) then
      if (row = char_rom_rows) then
        data <= (others => '0');
      else
        data <= read_data;
     end if;
    end if;
  end process;

end;

------------------------------- end of file --------------------------------
